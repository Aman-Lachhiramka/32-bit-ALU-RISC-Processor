`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.05.2023 14:01:05
// Design Name: 
// Module Name: adder_tb1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module alu_tb;
reg [31:0] x1;
reg [31:0] x2;
wire [31:0] x3;
reg [2:0] OpCode;
reg clk;

alu dut(.OpCode(OpCode),.x1(x1),.x2(x2),.x3(x3),.clk(clk));

always
#2 clk=~clk;

initial begin
clk=1;
OpCode = 3'b000;
x1= 32'b01000000010010010000111111011011;             //3.14
x2=32'b01000000100101010111000010100100    ;             //4.67


#5 
OpCode = 3'b001;
x1= 32'b01000000010010010000111111011011;             //3.14
x2=32'b01000000100101010111000010100100    ;             //4.67


#5
OpCode =3'b000;
x1= 32'b01000000010010001111010111000011;             //3.14
x2=32'b11000000010010001111010111000011    ;             //-3.14

#5
OpCode =3'b001;
x1= 32'b01000000010010001111010111000011;             //3.14
x2=32'b11000000010010001111010111000011    ;             //-3.14

//#5 x1= 32'b01000000010010010000111111011011;             //3.14
//x2=32'b11000000000100001010001111010111    ;             //-2.26

//#5 x1= 32'b11000000010010001111010111000011 ;             //-3.14
//x2=32'b11000000000100001010001111010111    ;             //-2.26

//#5 x1= 32'b11000001000101000010100011110110 ;             //-9.26
//x2=32'b11000000000100001010001111010111    ;             //-2.26

//#5 x1= 32'b01000001000101000010100011110110 ;             //9.26
//x2=32'b01000000000100001010001111010111    ;             //2.26

#5 
OpCode =3'b000;
x1= 32'b00000000000000000000000000000000 ;             //0
x2=32'b01111111100000000000000000000000    ;             //infinity

#5
OpCode =3'b000;
x1= 32'b01111111100000000000000000000000 ;             //infinity
x2=32'b01111111100000000000000000000000    ;             //infinity


// 45.13 * 63.13 = 2849.0569
#5
OpCode = 3'b011;
x1=32'h4234851F;
x2=32'h427C851F;

#5
//3.15 * -14.39 = -45.3285
x1=32'h4049999A;
x2=32'hC1663D71;

#5
//-13.15 * -48.16 = 633.304
x1=32'hC1526666;
x2=32'hC240A3D7;

#5
//inf*inf
x1=32'h7F800000;
x2=32'h7F800000;


#5
//-inf*inf
x1=32'b11111111100000000000000000000000;
x2=32'h7F800000;


#5
//-inf*-inf
x1=32'b11111111100000000000000000000000;
x2=32'b11111111100000000000000000000000;


//Testbench of OR
#5
OpCode=3'b101;
x1=32'b11111111100000000000000000000000;
x2=32'b11111111100000000000000000000000;

#5
x1=32'b11111111100000000000000111000000;
x2=32'b11111111100000000010000000000100;

//Testbench of AND
#5
OpCode=3'b100;
x1=32'b11111111100000000000000000000000;
x2=32'b11111111100000000000000000000000;

#5
x1=32'b11111111100000000000000111000000;
x2=32'b11111111100000000010000000000100;

//Testbench of XOR
#5
OpCode=3'b110;
x1=32'b11111111100000000000000000000000;
x2=32'b11111111100000000000000000000000;

#5
x1=32'b11111111100000000000000111000000;
x2=32'b11111111100000000010000000000100;


end
endmodule