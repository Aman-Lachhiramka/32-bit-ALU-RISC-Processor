`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.05.2023 16:42:29
// Design Name: 
// Module Name: adder_subtracter_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.05.2023 14:01:05
// Design Name: 
// Module Name: adder_tb1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module adder_subtracter_tb;
reg [31:0] x1;
reg [31:0] x2;
wire [31:0] x3;

adder_subtracter dut(.x1(x1),.x2(x2),.x3(x3));

initial begin
#5 x1= 32'b01000000010010010000111111011011;             //3.14
x2=32'b01000000100101010111000010100100    ;             //4.67

#5 x1= 32'b01000000010010001111010111000011;             //3.14
x2=32'b11000000010010001111010111000011    ;             //-3.14

#5 x1= 32'b01000000010010010000111111011011;             //3.14
x2=32'b11000000000100001010001111010111    ;             //-2.26

#5 x1= 32'b11000000010010001111010111000011 ;             //-3.14
x2=32'b11000000000100001010001111010111    ;             //-2.26

#5 x1= 32'b11000001000101000010100011110110 ;             //-9.26
x2=32'b11000000000100001010001111010111    ;             //-2.26

#5 x1= 32'b01000001000101000010100011110110 ;             //9.26
x2=32'b01000000000100001010001111010111    ;             //2.26

#5 x1= 32'b00000000000000000000000000000000 ;             //0
x2=32'b01111111100000000000000000000000    ;             //infinity

#5 x1= 32'b01111111100000000000000000000000 ;             //infinity
x2=32'b01111111100000000000000000000000    ;             //infinity

//#5 x1= 32'b01111111100000000000000000000001 ;             //NAN
//x2=32'b01111111100000000000000000000001   ;             //NAN

#5 x1= 32'b01111111100000000000000000000000 ;             //infinity
x2=32'b11111111100000000000000000000000    ;             //-infinity


////---
//#5 x1= 32'b01111111100000000000000000000001 ;             //NAN
//x2=32'b01000000000100001010001111010111   ;             //2.26

#5 x1= 32'b01111111100000000000000000000000 ;             //INFINITY
x2=32'b01000000000100001010001111010111   ;             //2.26

//#5 x1= 32'b01111111100000000000000000000000 ;             //infinity
//x2=32'b01111111100000000000000000000001   ;             //NAN

//#5 x1= 32'b01111111100000000000000000000001 ;             //NAN
//x2=32'b01111111100000000000000000000000  ;             //infi


end
endmodule
